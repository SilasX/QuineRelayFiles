module QR;initial begin $write("   \t\t\t \t\t\t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t \t\t\t\t\t\n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t \t\t\t\t\t\n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t \t    \n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t \t\t\t\t\t\n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t \t   \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("    \t \t   \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("    \t \t   \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("    \t \t   \n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("    \t \t   \n\t\n  ");$write("    \t \t   \n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t\t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("    \t \t   \n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("    \t \t   \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t\t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("    \t \t   \n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("    \t \t   \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t \t    \n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("    \t \t   \n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t \t   \n\t\n  ");$write("    \t \t   \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t \t   \n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("   \t \t\t\t \t\n\t\n  ");$write("    \t \t   \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t \t   \n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("    \t \t   \n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("    \t \t   \n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t\t\t\t \t \n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("    \t \t   \n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("    \t \t   \n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t     \n\t\n  ");$write("    \t     \n\t\n  ");$write("    \t     \n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t  \t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("    \t \t   \n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("    \t \t   \n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("    \t \t   \n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("   \t \t\t\t \t\n\t\n  ");$write("    \t \t   \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("    \t \t   \n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t \t   \n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("    \t \t   \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t \t   \n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("    \t \t   \n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("    \t \t   \n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("    \t \t   \n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t     \n\t\n  ");$write("    \t     \n\t\n  ");$write("    \t     \n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("   \t \t\t\t \t\n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("    \t \t   \n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("    \t \t   \n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("    \t     \n\t\n  ");$write("    \t   \t\t\n\t\n  ");$write("    \t \t   \n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("    \t \t   \n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t     \n\t\n  ");$write("    \t     \n\t\n  ");$write("    \t     \n\t\n  ");$write("    \t     \n\t\n  ");$write("    \t     \n\t\n  ");$write("    \t     \n\t\n  ");$write("    \t     \n\t\n  ");$write("    \t     \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t  \t \t\n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("    \t \t   \n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t\t\t\t \t \n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("   \t \t    \n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("   \t \t    \n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("   \t \t\t\t \t\n\t\n  ");$write("    \t \t   \n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("   \t \t    \n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t \t   \n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("    \t \t   \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t\t \t \t\t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("    \t \t   \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("    \t \t   \n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t \t    \n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("    \t \t   \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t \t   \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t  \t  \n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("    \t \t   \n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t \t   \n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("    \t   \t\t\n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("    \t \t   \n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("    \t     \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("    \t     \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t \t   \n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("    \t \t   \n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("    \t \t \t \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("    \t \t   \n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("    \t     \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t  \t  \n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t\t \t \t\t\n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t     \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t  \t  \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t \t   \n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("    \t     \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t  \t  \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("    \t \t   \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t     \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("   \t \t    \n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("   \t    \t \n\t\n  ");$write("    \t   \t\t\n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("    \t   \t\t\n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("    \t \t   \n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("    \t \t   \n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("    \t \t   \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("   \t \t\t\t \t\n\t\n  ");$write("   \t \t\t\t\t\t\n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t \t\t\t\t\t\n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("   \t \t    \n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t \t    \n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("   \t \t    \n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("    \t \t   \n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("    \t \t   \n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t\t \t \t\t\n\t\n  ");$write("    \t     \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("   \t \t    \n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("    \t \t   \n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("   \t \t\t\t \t\n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("   \t \t\t\t \t\n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t \t\t\t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t\t\t\t \t \n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t    \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t \t\t\n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t     \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t    \t \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t    \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t    \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t\t\t\t \t \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t \t    \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t    \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t\t \t \t\t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t     \t\n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t \t    \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t    \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t    \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t\t\t\t \t \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("   \t\t \t \t\t\n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("   \t\t\t\t \t \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t\t \t \t\t\n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t\t\t\t \t \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("   \t    \t \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t    \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("   \t \t    \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t    \t \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t    \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t    \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t    \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t \t    \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t \t \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t    \t \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("   \t\t \t \t\t\n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t\t\t\t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t\t \t \t\t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t \t    \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t     \t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t\t \t \t\t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t     \t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t \t    \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t    \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t\t\t \t \n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t     \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("   \t\t\t\t \t \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("   \t     \t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t     \t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t \t \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t \t \t\t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("   \t \t    \n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t\t \t \t\t\n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("   \t\t \t \t\t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t\t\t\t \t \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("   \t \t    \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("   \t\t \t \t\t\n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("   \t     \t\n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("   \t    \t \n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("   \t    \t \n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t    \t \n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t\t\t\t \t \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("   \t    \t \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("   \t\t \t \t\t\n\t\n  ");$write("   \t    \t \n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("   \t    \t \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t \t    \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t\t \t \t\t\n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t\t \t \t\t\n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t    \n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("   \t    \t \n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("   \t    \t \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("   \t\t \t \t\t\n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("   \t    \t \n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t    \t \n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("   \t    \t \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("   \t    \t \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t    \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t \t    \n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("   \t\t\t\t \t \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("   \t \t    \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("   \t \t    \n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("   \t\t \t \t\t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t\t \t \t\t\n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("   \t    \t \n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("   \t    \t \n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t \t \n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("   \t\t\t\t \t \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("   \t     \t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t    \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("   \t\t\t\t \t \n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("   \t \t    \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("   \t \t    \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("   \t\t \t \t\t\n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t\t\t\t \t \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t    \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t \t    \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("   \t\t \t \t\t\n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t \t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t    \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t\t\t\t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t    \n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("   \t    \t \n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("   \t    \t \n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("   \t    \t \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t    \t \n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t    \t \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t     \t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t    \t \n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t\t\t\t \t \n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t \t    \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("   \t \t    \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t\t \t \t\t\n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("   \t \t    \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t     \t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("   \t \t    \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("   \t \t    \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t    \t \n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t    \n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("   \t \t    \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t \t    \n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t    \n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("   \t     \t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t    \t \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("   \t \t    \n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t \t    \n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("   \t \t    \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t\t\t\t \t \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("   \t    \t \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("   \t    \t \n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("   \t \t    \n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("   \t \t    \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("   \t \t    \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t \t    \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t \t    \n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("   \t \t    \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t\t\t\t \t \n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t \t    \n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t    \t \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("   \t\t \t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("   \t\t \t \t\t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("   \t \t    \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t \t    \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t    \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t    \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("   \t    \t \n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t\t \t \t\t\n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("   \t \t    \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t \t    \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("   \t    \t \n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("   \t \t    \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("   \t \t    \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t \t    \n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("   \t\t\t\t \t \n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("   \t \t    \n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("   \t    \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("   \t    \t \n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t\t \t \t\t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("   \t\t \t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("   \t \t    \n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t \t    \n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("   \t \t    \n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t \t    \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("   \t \t    \n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("   \t\t\t\t \t \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("   \t\t\t\t \t \n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("   \t \t    \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("   \t \t    \n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("   \t    \t \n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t\t \t \t\t\n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t    \n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("   \t    \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t \t \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t \t    \n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t    \n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t\t \t \t\t\n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("   \t \t    \n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("   \t \t    \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("   \t\t \t \t\t\n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t \t    \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("   \t\t \t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("   \t\t \t \t\t\n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t \t    \n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("   \t\t \t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t\t \t \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t    \t \n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("   \t    \t \n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("   \t    \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t \t \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t    \t \n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t \t \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t \t    \n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("   \t    \t \n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("   \t\t\t\t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t    \t \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("   \t    \t \n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("   \t \t    \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t\t\t\t \t \n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("   \t    \t \n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("   \t\t\t\t \t \n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("   \t\t \t \t\t\n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t \t    \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t \t    \n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t     \t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t \t    \n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t    \t \n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t    \t \n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t    \n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t \t    \n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("   \t \t    \n\t\n  ");$write("   \t\t \t \t\t\n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t    \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("   \t \t    \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("   \t \t    \n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("   \t\t\t\t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("   \t \t    \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("   \t \t    \n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("   \t\t\t\t \t \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("   \t\t\t\t \t \n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("   \t \t    \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t    \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t    \n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t    \t \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("   \t    \t \n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("   \t \t    \n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("   \t\t\t\t \t \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("   \t\t \t \t\t\n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t    \t \n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t    \t \n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("   \t\t \t \t\t\n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("   \t \t    \n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("   \t \t    \n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("   \t    \t \n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t \t    \n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t \t    \n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("   \t\t \t \t\t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("   \t     \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("   \t \t    \n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("   \t\t \t \t\t\n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("   \t\t \t \t\t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("   \t \t    \n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("   \t \t    \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("   \t \t    \n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("   \t\t \t \t\t\n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("   \t \t    \n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("   \t\t \t \t\t\n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t \t    \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("   \t \t    \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t\t \t \t\t\n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t \t    \n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t \t \n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("   \t\t \t \t\t\n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t \t    \n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("   \t\t\t\t \t \n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t\t\t\t \t \n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t \t \t\t\n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t    \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("   \t \t    \n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("   \t\t\t\t \t \n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("   \t\t \t \t\t\n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t \t    \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t \t    \n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("   \t    \t \n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("   \t\t \t \t\t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("   \t\t \t \t\t\n\t\n  ");$write("   \t\t \t \t\t\n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("   \t \t    \n\t\n  ");$write("   \t\t \t \t\t\n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t    \t \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("   \t\t\t\t \t \n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t \t    \n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("   \t\t\t\t \t \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("   \t\t \t \t\t\n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("   \t\t\t\t \t \n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t    \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t \t    \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t\t \t \t\t\n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("   \t\t \t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t\t \t \t\t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("   \t \t    \n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("   \t \t    \n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("   \t\t \t \t\t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t \t \n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t\t \t \t\t\n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("   \t\t\t\t \t \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t \t    \n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t    \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t \t    \n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("   \t\t \t \t\t\n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t    \n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("   \t \t    \n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t\t\t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t \t    \n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("   \t\t \t \t\t\n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("   \t\t\t\t \t \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("   \t\t \t \t\t\n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("   \t \t    \n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("   \t\t \t \t\t\n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t\t \t \t\t\n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("   \t    \t \n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("   \t\t\t\t \t \n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t\t \t \t\t\n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("   \t \t    \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("   \t\t\t\t \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("   \t\t \t \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t\t \t \t\t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("   \t\t \t \t\t\n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t\t \t \t\t\n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t\t\t\t \t \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("   \t\t\t\t \t \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("   \t \t    \n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t    \n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("   \t\t \t \t\t\n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t\t \t \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("   \t\t \t \t\t\n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t\t \t \t\t\n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("   \t\t \t \t\t\n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("   \t\t \t \t\t\n\t\n  ");$write("   \t \t    \n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("   \t\t \t \t\t\n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("   \t\t\t\t \t \n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t    \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("   \t\t \t \t\t\n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("   \t \t    \n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("   \t\t\t\t \t \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("   \t \t    \n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("   \t     \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t\t \t \t\t\n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("   \t\t \t \t\t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("   \t\t \t \t\t\n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t    \n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("   \t\t\t\t \t \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("   \t\t\t\t \t \n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("   \t    \t \n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("   \t \t    \n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t \t \n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("   \t\t \t \t\t\n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t\t\t\t \t \n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("   \t    \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("   \t\t \t \t\t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("   \t     \t\n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("   \t \t    \n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t\t \t \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t \t \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t\t \t \t\t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("   \t\t \t \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("   \t    \t \n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("   \t \t    \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t\t\t\t \t \n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t \t    \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t \t    \n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t \t    \n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t    \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("   \t \t    \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("   \t    \t \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("   \t\t\t\t \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t \t    \n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t \t    \n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("   \t \t    \n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t \t    \n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t  \t\t \t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t     \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t    \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("   \t  \t   \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t    \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("   \t\t \t \t\t\n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t \t\t\n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t\t \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("   \t \t    \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t  \t \t\t\n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t \t    \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("    \t\t\t   \n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t\t\t\t \t \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t \t\t   \n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("    \t \t   \n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t \t\t\t \t\n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("    \t \t   \n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("    \t \t   \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("    \t \t   \n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("    \t \t   \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("    \t \t \t \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("    \t\t \t\t \n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("    \t\t\t  \t\n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("    \t \t \t \n\t\n  ");$write("    \t\t \t \t\n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("    \t\t \t  \n\t\n  ");$write("    \t\t  \t\t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t \t   \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t  \t \t\n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("   \t\t\t\t \t\t\n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("    \t\t\t\t\t\t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("   \t \t\t\t \t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t \t\t\t \t\n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("   \t\t\t\t \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("    \t \t   \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("    \t \t   \n\t\n  ");$write("   \t\t\t\t \t \n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("   \t \t\t\t \t\n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t\t   \t\n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t\t\t\t \t\n\t\n  ");$write("   \t\t\t\t\t \t\n\t\n  ");$write("   \t\t\t\t\t \t\n\t\n  ");$write("   \t\t\t\t\t \t\n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("   \t\t \t \t\t\n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("   \t \t    \n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("    \t \t   \n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t\t\t \t\t \n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("   \t \t \t\t \n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("    \t\t  \t \n\t\n  ");$write("    \t\t \t\t\t\n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("   \t      \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("    \t\t   \t\n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("   \t\t\t\t\t \t\n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t     \n\t\n  ");$write("    \t     \n\t\n  ");$write("    \t     \n\t\n  ");$write("    \t     \n\t\n  ");$write("    \t     \n\t\n  ");$write("    \t     \n\t\n  ");$write("    \t     \n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("    \t \t   \n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t     \n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("   \t \t\t\t \t\n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t   \n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t   \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("    \t \t   \n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("   \t \t    \n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t \t   \n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("    \t \t   \n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t \t   \n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("    \t \t   \n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("    \t \t   \n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("   \t \t    \n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t \t   \n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("    \t \t   \n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("    \t \t   \n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("    \t \t   \n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("   \t \t    \n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t \t   \n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("    \t \t   \n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("    \t \t\t \t\n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("   \t \t \t\t\t\n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("    \t \t   \n\t\n  ");$write("    \t \t \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t \t \t \n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("    \t  \t\t\t\n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t  \t\t\t\n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("    \t \t   \n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("   \t \t    \n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t \t   \n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t \t   \n\t\n  ");$write("    \t  \t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("    \t \t   \n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("   \t \t    \n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t \t   \n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t  \t\t \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t  \t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("    \t \t   \n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("   \t \t    \n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t \t   \n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t  \t\t \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t  \t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t\t\t\t \t\n\t\n  ");$write("    \t\t    \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("    \t \t   \n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("   \t \t    \n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t \t   \n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t  \t\t \n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("    \t \t   \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("   \t    \t\t\n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("    \t \t   \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t  \t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("   \t\t\t \t\t\t\n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t\t\t\t  \n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t\t \t   \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("    \t \t   \n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t  \t  \t\n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("   \t \t    \n\t\n  ");$write("   \t  \t\t  \n\t\n  ");$write("   \t     \t\n\t\n  ");$write("   \t \t\t  \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t \t   \n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t  \t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t\t \t\t \t\n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("   \t \t    \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("   \t\t\t\t  \t\n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("   \t \t  \t\t\n\t\n  ");$write("   \t \t \t  \n\t\n  ");$write("   \t  \t\t\t\t\n\t\n  ");$write("   \t \t    \n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("   \t \t \t \t\n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("   \t \t\t\t \t\n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("   \t\t \t\t  \n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t\t   \t\t\n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t \t   \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("   \t\t\t\t\t\t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t\t\t\t \t\n\t\n  ");$write("   \t\t\t\t\t \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t\t\t\t \t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("    \t     \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t\t\t\t \t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("    \t\t\t \t \n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t\t \t \t \n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("    \t \t   \n\t\n  ");$write("   \t \t\t \t\t\n\t\n  ");$write("    \t  \t\t\t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("    \t  \t\t\t\n\t\n  ");$write("   \t\t  \t\t \n\t\n  ");$write("   \t\t \t\t\t\t\n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("   \t\t    \t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("    \t \t   \n\t\n  ");$write("    \t\t    \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("   \t \t\t\t \t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("    \t \t \t\t\n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t \t\t\t \n\t\n  ");$write("    \t\t\t\t\t \n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t  \t\t\t\n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("   \t\t\t \t \t\n\t\n  ");$write("   \t\t   \t \n\t\n  ");$write("    \t \t   \n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("    \t    \t\n\t\n  ");$write("    \t \t\t\t\t\n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("   \t \t\t\t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t \t\t  \n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t\t    \n\t\n  ");$write("   \t\t\t  \t \n\t\n  ");$write("   \t\t \t  \t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t\t\t \t  \n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t\t\t  \t\t\n\t\n  ");$write("   \t\t\t\t\t \t\n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("   \t   \t \t\n\t\n  ");$write("   \t  \t\t\t \n\t\n  ");$write("   \t   \t  \n\t\n  ");$write("    \t   \t \n\t\n  ");$write("    \t \t  \t\n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$write("   \t\t  \t \t\n\t\n  ");$write("   \t\t \t\t\t \n\t\n  ");$write("   \t\t  \t  \n\t\n  ");$write("    \t     \n\t\n  ");$write("   \t \t   \t\n\t\n  ");$write("   \t \t  \t \n\t\n  ");$write("    \t\t\t \t\t\n\t\n  ");$display("\n\n");end endmodule